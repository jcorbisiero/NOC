module noc
(
	ifc.nic n
);




endmodule


