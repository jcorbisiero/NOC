module noc
(
	ifc_noc.noc n
);




endmodule


